module judge(

   );
endmodule